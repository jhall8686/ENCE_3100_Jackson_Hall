module seg_decoder(
	input[2:0] c,
	output[7:0] m
	);
	wire m12;
	mux_2_1(c[2], ~(c[2] | c[0]), 1, m[0]);
	mux_2_1(c[2], (c[1] ^ c[0]), 1, m12);
	assign m12 = m[1];
	assign m12 = m[2];
	mux_2_1(c[2], ~(c[1] | c[0]), 1, m[3]);
	assign m[4] = c[2];
	assign m[5] = c[2];
	mux_2_1(c[2], (c[1] & ~c[0]), 1, m[6]);
	assign m[7] = 1;
	
endmodule
	