module BCD_decoder(
	input [3:0] bcd,
	output [7:0] seg
	);
	
	always @(*) begin
		case(bcd)
			4'd0: 8'b00000011;
			4'd1:	8'b10011111;
			4'd2:	8'b00100101;
			4'd3:	8'b00001101;
			4'd4: 8'b10011001;
			4'd5: 8'b01001001;
			4'd6:	8'b01000001;
			4'd7: 8'b00011111;
			4'd8: 8'b00000001;
			4'd9: 8'b00001001;
			4'd10: 8'b11111111;
			4'd11: 8'b11111111;
			4'd12: 8'b11111111;
			4'd13: 8'b11111111;
			4'd14: 8'b11111111;
			4'd15: 8'b11111111;
			default:
		endcase
	end
	
	
	
endmodule